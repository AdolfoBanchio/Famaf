module maindec(input logic [10:0]op,
					input logic reset,
					output logic Reg2Loc,MemtoReg,RegWrite,
					MemRead,MemWrite,Branch,NotAnInstr,ERet,
					output logic [1:0]ALUOp,ALUSrc);
	always_comb begin
		if (!reset) begin
			casez(op)
			//R-format
				'b100_0101_1000:begin
								Reg2Loc='b0;
								ALUSrc='b00;
								MemtoReg='b0;
								RegWrite='b1;
								MemRead='b0;
								MemWrite='b0;
								Branch='b0;
								ALUOp='b10;
								NotAnInstr='b0;
								ERet='b0;
								end
				'b110_0101_1000:begin
								Reg2Loc='b0;
								ALUSrc='b00;
								MemtoReg='b0;
								RegWrite='b1;
								MemRead='b0;
								MemWrite='b0;
								Branch='b0;
								ALUOp='b10;
								NotAnInstr='b0;
								ERet='b0;
								end
				'b100_0101_0000:begin
								Reg2Loc='b0;
								ALUSrc='b00;
								MemtoReg='b0;
								RegWrite='b1;
								MemRead='b0;
								MemWrite='b0;
								Branch='b0;
								ALUOp='b10;
								NotAnInstr='b0;
								ERet='b0;
								end
				'b101_0101_0000:begin
								Reg2Loc='b0;
								ALUSrc='b00;
								MemtoReg='b0;
								RegWrite='b1;
								MemRead='b0;
								MemWrite='b0;
								Branch='b0;
								ALUOp='b10;
								NotAnInstr='b0;
								ERet='b0;
								end
                 //BR
				'b110_1011_0000:begin
								Reg2Loc='b0;
								ALUSrc='b00;
								MemtoReg='b0;
								RegWrite='b0;
								MemRead='b0;
								MemWrite='b0;
								Branch='b0;
								ALUOp='b10;
								NotAnInstr='b0;
								ERet='b0;
								end
				//ERET
				'b1101011_0100:begin
								Reg2Loc='b0;
								ALUSrc='b00;
								MemtoReg='bX;
								RegWrite='b0;
								MemRead='b0;
								MemWrite='b0;
								Branch='b1;
								ALUOp='b01;
								NotAnInstr='b0;
								ERet='b1;
								end
				//MRS
				'b110_1010_1001:begin
								Reg2Loc='b1;
								ALUSrc='b1X;
								MemtoReg='b0;
								RegWrite='b1;
								MemRead='b0;
								MemWrite='b0;
								Branch='b0;
								ALUOp='b01;
								NotAnInstr='b0;
								ERet='b0;
								end
				//LDUR
				'b111_1100_0010:begin
								Reg2Loc='b0;
								ALUSrc='b01;
								MemtoReg='b1;
								RegWrite='b1;
								MemRead='b1;
								MemWrite='b0;
								Branch='b0;
								ALUOp='b00;
								NotAnInstr='b0;
								ERet='b0;
								end
				//STUR
				'b111_1100_0000:begin
								Reg2Loc='b1;
								ALUSrc='b01;
								MemtoReg='b0;
								RegWrite='b0;
								MemRead='b0;
								MemWrite='b1;
								Branch='b0;
								ALUOp='b00;
								NotAnInstr='b0;
								ERet='b0;
								end
				//CBZ
				'b101_1010_0???:begin
								Reg2Loc='b1;
								ALUSrc='b00;
								MemtoReg='b0;
								RegWrite='b0;
								MemRead='b0;
								MemWrite='b0;
								Branch='b1;
								ALUOp='b01;
								NotAnInstr='b0;
								ERet='b0;
								end
				default: begin
						 Reg2Loc='bX;
						 ALUSrc='bXX;
						 MemtoReg='b0;
						 RegWrite='b0;
						 MemRead='b0;
						 MemWrite='b0;
						 Branch='b1;
						 ALUOp='bXX;
						 NotAnInstr='b1;
						 ERet='b0;
						 end
			endcase
		end else begin 
			Reg2Loc='b0;
			ALUSrc='b00;
			MemtoReg='b0;
			RegWrite='b0;
			MemRead='b0;
			MemWrite='b0;
			Branch='b0;
			ALUOp='b00;
			NotAnInstr='b0;
			ERet='b0;
		end
	end
endmodule