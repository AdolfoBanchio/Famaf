module maindec(input logic [10:0]op,
			   output logic Reg2Loc,ALUSrc,MemtoReg,RegWrite,
			   MemRead,MemWrite,Branch,
			   output logic [1:0]ALUOp);
	always_comb begin
		casez(op)
		//R-format
			'b100_0101_1000:begin
							Reg2Loc='b0;
							ALUSrc='b0;
							MemtoReg='b0;
							RegWrite='b1;
							MemRead='b0;
							MemWrite='b0;
							Branch='b0;
							ALUOp='b10;
							end
			'b110_0101_1000:begin
							Reg2Loc='b0;
							ALUSrc='b0;
							MemtoReg='b0;
							RegWrite='b1;
							MemRead='b0;
							MemWrite='b0;
							Branch='b0;
							ALUOp='b10;
							end
			'b100_0101_0000:begin
							Reg2Loc='b0;
							ALUSrc='b0;
							MemtoReg='b0;
							RegWrite='b1;
							MemRead='b0;
							MemWrite='b0;
							Branch='b0;
							ALUOp='b10;
							end
			'b101_0101_0000:begin
							Reg2Loc='b0;
							ALUSrc='b0;
							MemtoReg='b0;
							RegWrite='b1;
							MemRead='b0;
							MemWrite='b0;
							Branch='b0;
							ALUOp='b10;
							end
			//LDUR
			'b111_1100_0010:begin
							Reg2Loc='b0;
							ALUSrc='b1;
							MemtoReg='b1;
							RegWrite='b1;
							MemRead='b1;
							MemWrite='b0;
							Branch='b0;
							ALUOp='b00;
							end
			//STUR
			'b111_1100_0000:begin
							Reg2Loc='b1;
							ALUSrc='b1;
							MemtoReg='b0;
							RegWrite='b0;
							MemRead='b0;
							MemWrite='b1;
							Branch='b0;
							ALUOp='b00;
							end
			//CBZ
			'b101_1010_0???:begin
							Reg2Loc='b1;
							ALUSrc='b0;
							MemtoReg='b0;
							RegWrite='b0;
							MemRead='b0;
							MemWrite='b0;
							Branch='b1;
							ALUOp='b01;
							end
			default: begin
					 Reg2Loc='b1;
					 ALUSrc='b0;
					 MemtoReg='b0;
					 RegWrite='b0;
					 MemRead='b0;
					 MemWrite='b0;
					 Branch='b1;
					 ALUOp='b01;
					 end
		endcase
	end
endmodule